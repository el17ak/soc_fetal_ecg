// Computer_System.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module Computer_System (
		input  wire [31:0] hps_f2h_irq0_irq,                //         hps_f2h_irq0.irq
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                     .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                     .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                     .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                     .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                     .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                     .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //                     .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                     .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                    //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                     .mem_ba
		output wire        memory_mem_ck,                   //                     .mem_ck
		output wire        memory_mem_ck_n,                 //                     .mem_ck_n
		output wire        memory_mem_cke,                  //                     .mem_cke
		output wire        memory_mem_cs_n,                 //                     .mem_cs_n
		output wire        memory_mem_ras_n,                //                     .mem_ras_n
		output wire        memory_mem_cas_n,                //                     .mem_cas_n
		output wire        memory_mem_we_n,                 //                     .mem_we_n
		output wire        memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire        memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                     .mem_dm
		input  wire        memory_oct_rzqin,                //                     .oct_rzqin
		input  wire        onchip_sram_clk2_clk,            //     onchip_sram_clk2.clk
		input  wire        onchip_sram_reset2_reset,        //   onchip_sram_reset2.reset
		input  wire        onchip_sram_reset2_reset_req,    //                     .reset_req
		input  wire [13:0] onchip_sram_s2_address,          //       onchip_sram_s2.address
		input  wire        onchip_sram_s2_chipselect,       //                     .chipselect
		input  wire        onchip_sram_s2_clken,            //                     .clken
		input  wire        onchip_sram_s2_write,            //                     .write
		output wire [31:0] onchip_sram_s2_readdata,         //                     .readdata
		input  wire [31:0] onchip_sram_s2_writedata,        //                     .writedata
		input  wire [3:0]  onchip_sram_s2_byteenable,       //                     .byteenable
		output wire        sdram_clk_clk,                   //            sdram_clk.clk
		input  wire        system_pll_ref_clk_clk,          //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset       // system_pll_ref_reset.reset
	);

	wire         system_pll_sys_clk_clk;                                // System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, Onchip_SRAM:clk, dma_1:clk, dma_2:clk, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, mm_interconnect_2:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk]
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                  // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                    // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                    // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire         arm_a9_hps_h2f_lw_axi_master_wready;                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                      // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire         arm_a9_hps_h2f_lw_axi_master_rready;                   // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                    // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                      // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                  // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire         arm_a9_hps_h2f_lw_axi_master_wvalid;                   // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                   // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                   // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                   // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                    // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire         arm_a9_hps_h2f_lw_axi_master_arvalid;                  // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                  // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                     // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                   // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                   // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                   // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire         arm_a9_hps_h2f_lw_axi_master_arready;                  // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire         arm_a9_hps_h2f_lw_axi_master_awready;                  // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                  // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                   // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire         arm_a9_hps_h2f_lw_axi_master_bready;                   // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire         arm_a9_hps_h2f_lw_axi_master_rlast;                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire         arm_a9_hps_h2f_lw_axi_master_wlast;                    // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                    // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                     // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                      // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire         arm_a9_hps_h2f_lw_axi_master_bvalid;                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                   // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire         arm_a9_hps_h2f_lw_axi_master_awvalid;                  // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire         arm_a9_hps_h2f_lw_axi_master_rvalid;                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire         mm_interconnect_0_dma_1_control_port_slave_chipselect; // mm_interconnect_0:dma_1_control_port_slave_chipselect -> dma_1:dma_ctl_chipselect
	wire  [31:0] mm_interconnect_0_dma_1_control_port_slave_readdata;   // dma_1:dma_ctl_readdata -> mm_interconnect_0:dma_1_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_1_control_port_slave_address;    // mm_interconnect_0:dma_1_control_port_slave_address -> dma_1:dma_ctl_address
	wire         mm_interconnect_0_dma_1_control_port_slave_write;      // mm_interconnect_0:dma_1_control_port_slave_write -> dma_1:dma_ctl_write_n
	wire  [31:0] mm_interconnect_0_dma_1_control_port_slave_writedata;  // mm_interconnect_0:dma_1_control_port_slave_writedata -> dma_1:dma_ctl_writedata
	wire         mm_interconnect_0_dma_2_control_port_slave_chipselect; // mm_interconnect_0:dma_2_control_port_slave_chipselect -> dma_2:dma_ctl_chipselect
	wire  [31:0] mm_interconnect_0_dma_2_control_port_slave_readdata;   // dma_2:dma_ctl_readdata -> mm_interconnect_0:dma_2_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_2_control_port_slave_address;    // mm_interconnect_0:dma_2_control_port_slave_address -> dma_2:dma_ctl_address
	wire         mm_interconnect_0_dma_2_control_port_slave_write;      // mm_interconnect_0:dma_2_control_port_slave_write -> dma_2:dma_ctl_write_n
	wire  [31:0] mm_interconnect_0_dma_2_control_port_slave_writedata;  // mm_interconnect_0:dma_2_control_port_slave_writedata -> dma_2:dma_ctl_writedata
	wire         dma_1_read_master_chipselect;                          // dma_1:read_chipselect -> mm_interconnect_1:dma_1_read_master_chipselect
	wire  [31:0] dma_1_read_master_readdata;                            // mm_interconnect_1:dma_1_read_master_readdata -> dma_1:read_readdata
	wire         dma_1_read_master_waitrequest;                         // mm_interconnect_1:dma_1_read_master_waitrequest -> dma_1:read_waitrequest
	wire  [31:0] dma_1_read_master_address;                             // dma_1:read_address -> mm_interconnect_1:dma_1_read_master_address
	wire         dma_1_read_master_read;                                // dma_1:read_read_n -> mm_interconnect_1:dma_1_read_master_read
	wire         dma_1_read_master_readdatavalid;                       // mm_interconnect_1:dma_1_read_master_readdatavalid -> dma_1:read_readdatavalid
	wire         dma_2_write_master_chipselect;                         // dma_2:write_chipselect -> mm_interconnect_1:dma_2_write_master_chipselect
	wire         dma_2_write_master_waitrequest;                        // mm_interconnect_1:dma_2_write_master_waitrequest -> dma_2:write_waitrequest
	wire  [31:0] dma_2_write_master_address;                            // dma_2:write_address -> mm_interconnect_1:dma_2_write_master_address
	wire   [3:0] dma_2_write_master_byteenable;                         // dma_2:write_byteenable -> mm_interconnect_1:dma_2_write_master_byteenable
	wire         dma_2_write_master_write;                              // dma_2:write_write_n -> mm_interconnect_1:dma_2_write_master_write
	wire  [31:0] dma_2_write_master_writedata;                          // dma_2:write_writedata -> mm_interconnect_1:dma_2_write_master_writedata
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst;    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awburst -> ARM_A9_HPS:f2h_AWBURST
	wire   [4:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awuser -> ARM_A9_HPS:f2h_AWUSER
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen;      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlen -> ARM_A9_HPS:f2h_ARLEN
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb;      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wstrb -> ARM_A9_HPS:f2h_WSTRB
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready;     // ARM_A9_HPS:f2h_WREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid;        // ARM_A9_HPS:f2h_RID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rid
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rready -> ARM_A9_HPS:f2h_RREADY
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen;      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlen -> ARM_A9_HPS:f2h_AWLEN
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid;        // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wid -> ARM_A9_HPS:f2h_WID
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache;    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arcache -> ARM_A9_HPS:f2h_ARCACHE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wvalid -> ARM_A9_HPS:f2h_WVALID
	wire  [31:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_araddr -> ARM_A9_HPS:f2h_ARADDR
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arprot -> ARM_A9_HPS:f2h_ARPROT
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awprot -> ARM_A9_HPS:f2h_AWPROT
	wire  [63:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata;      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wdata -> ARM_A9_HPS:f2h_WDATA
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid;    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arvalid -> ARM_A9_HPS:f2h_ARVALID
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache;    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awcache -> ARM_A9_HPS:f2h_AWCACHE
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid;       // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arid -> ARM_A9_HPS:f2h_ARID
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlock -> ARM_A9_HPS:f2h_ARLOCK
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlock -> ARM_A9_HPS:f2h_AWLOCK
	wire  [31:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awaddr -> ARM_A9_HPS:f2h_AWADDR
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp;      // ARM_A9_HPS:f2h_BRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bresp
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready;    // ARM_A9_HPS:f2h_ARREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata;      // ARM_A9_HPS:f2h_RDATA -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rdata
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready;    // ARM_A9_HPS:f2h_AWREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst;    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arburst -> ARM_A9_HPS:f2h_ARBURST
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arsize -> ARM_A9_HPS:f2h_ARSIZE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bready -> ARM_A9_HPS:f2h_BREADY
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast;      // ARM_A9_HPS:f2h_RLAST -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rlast
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast;      // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wlast -> ARM_A9_HPS:f2h_WLAST
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp;      // ARM_A9_HPS:f2h_RRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid;       // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awid -> ARM_A9_HPS:f2h_AWID
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid;        // ARM_A9_HPS:f2h_BID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bid
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid;     // ARM_A9_HPS:f2h_BVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awsize -> ARM_A9_HPS:f2h_AWSIZE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid;    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awvalid -> ARM_A9_HPS:f2h_AWVALID
	wire   [4:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser;     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_aruser -> ARM_A9_HPS:f2h_ARUSER
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid;     // ARM_A9_HPS:f2h_RVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rvalid
	wire         dma_2_read_master_chipselect;                          // dma_2:read_chipselect -> mm_interconnect_2:dma_2_read_master_chipselect
	wire  [31:0] dma_2_read_master_readdata;                            // mm_interconnect_2:dma_2_read_master_readdata -> dma_2:read_readdata
	wire         dma_2_read_master_waitrequest;                         // mm_interconnect_2:dma_2_read_master_waitrequest -> dma_2:read_waitrequest
	wire  [27:0] dma_2_read_master_address;                             // dma_2:read_address -> mm_interconnect_2:dma_2_read_master_address
	wire         dma_2_read_master_read;                                // dma_2:read_read_n -> mm_interconnect_2:dma_2_read_master_read
	wire         dma_2_read_master_readdatavalid;                       // mm_interconnect_2:dma_2_read_master_readdatavalid -> dma_2:read_readdatavalid
	wire         dma_1_write_master_chipselect;                         // dma_1:write_chipselect -> mm_interconnect_2:dma_1_write_master_chipselect
	wire         dma_1_write_master_waitrequest;                        // mm_interconnect_2:dma_1_write_master_waitrequest -> dma_1:write_waitrequest
	wire  [27:0] dma_1_write_master_address;                            // dma_1:write_address -> mm_interconnect_2:dma_1_write_master_address
	wire   [3:0] dma_1_write_master_byteenable;                         // dma_1:write_byteenable -> mm_interconnect_2:dma_1_write_master_byteenable
	wire         dma_1_write_master_write;                              // dma_1:write_write_n -> mm_interconnect_2:dma_1_write_master_write
	wire  [31:0] dma_1_write_master_writedata;                          // dma_1:write_writedata -> mm_interconnect_2:dma_1_write_master_writedata
	wire         mm_interconnect_2_onchip_sram_s1_chipselect;           // mm_interconnect_2:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	wire  [31:0] mm_interconnect_2_onchip_sram_s1_readdata;             // Onchip_SRAM:readdata -> mm_interconnect_2:Onchip_SRAM_s1_readdata
	wire  [13:0] mm_interconnect_2_onchip_sram_s1_address;              // mm_interconnect_2:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	wire   [3:0] mm_interconnect_2_onchip_sram_s1_byteenable;           // mm_interconnect_2:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	wire         mm_interconnect_2_onchip_sram_s1_write;                // mm_interconnect_2:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	wire  [31:0] mm_interconnect_2_onchip_sram_s1_writedata;            // mm_interconnect_2:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	wire         mm_interconnect_2_onchip_sram_s1_clken;                // mm_interconnect_2:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;                               // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [Onchip_SRAM:reset, dma_1:system_reset_n, dma_2:system_reset_n, mm_interconnect_0:dma_1_reset_reset_bridge_in_reset_reset, mm_interconnect_1:dma_1_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	wire         arm_a9_hps_h2f_reset_reset;                            // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         system_pll_reset_source_reset;                         // System_PLL:reset_source_reset -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                                       //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                      //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                      //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                    //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                     //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                    //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                   //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                   //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                    //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                 //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                      //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                     //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                   //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                     //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                      //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                   //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                      //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                        //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                        //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                        //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                        //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                        //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                        //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),                     //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),                         //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                                   //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                                   //                  .awaddr
		.h2f_AWLEN                (),                                                   //                  .awlen
		.h2f_AWSIZE               (),                                                   //                  .awsize
		.h2f_AWBURST              (),                                                   //                  .awburst
		.h2f_AWLOCK               (),                                                   //                  .awlock
		.h2f_AWCACHE              (),                                                   //                  .awcache
		.h2f_AWPROT               (),                                                   //                  .awprot
		.h2f_AWVALID              (),                                                   //                  .awvalid
		.h2f_AWREADY              (),                                                   //                  .awready
		.h2f_WID                  (),                                                   //                  .wid
		.h2f_WDATA                (),                                                   //                  .wdata
		.h2f_WSTRB                (),                                                   //                  .wstrb
		.h2f_WLAST                (),                                                   //                  .wlast
		.h2f_WVALID               (),                                                   //                  .wvalid
		.h2f_WREADY               (),                                                   //                  .wready
		.h2f_BID                  (),                                                   //                  .bid
		.h2f_BRESP                (),                                                   //                  .bresp
		.h2f_BVALID               (),                                                   //                  .bvalid
		.h2f_BREADY               (),                                                   //                  .bready
		.h2f_ARID                 (),                                                   //                  .arid
		.h2f_ARADDR               (),                                                   //                  .araddr
		.h2f_ARLEN                (),                                                   //                  .arlen
		.h2f_ARSIZE               (),                                                   //                  .arsize
		.h2f_ARBURST              (),                                                   //                  .arburst
		.h2f_ARLOCK               (),                                                   //                  .arlock
		.h2f_ARCACHE              (),                                                   //                  .arcache
		.h2f_ARPROT               (),                                                   //                  .arprot
		.h2f_ARVALID              (),                                                   //                  .arvalid
		.h2f_ARREADY              (),                                                   //                  .arready
		.h2f_RID                  (),                                                   //                  .rid
		.h2f_RDATA                (),                                                   //                  .rdata
		.h2f_RRESP                (),                                                   //                  .rresp
		.h2f_RLAST                (),                                                   //                  .rlast
		.h2f_RVALID               (),                                                   //                  .rvalid
		.h2f_RREADY               (),                                                   //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0               (hps_f2h_irq0_irq),                                   //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	Computer_System_Onchip_SRAM onchip_sram (
		.clk         (system_pll_sys_clk_clk),                      //   clk1.clk
		.address     (mm_interconnect_2_onchip_sram_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_onchip_sram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_onchip_sram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_onchip_sram_s1_write),      //       .write
		.readdata    (mm_interconnect_2_onchip_sram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_onchip_sram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_onchip_sram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (onchip_sram_s2_address),                      //     s2.address
		.chipselect2 (onchip_sram_s2_chipselect),                   //       .chipselect
		.clken2      (onchip_sram_s2_clken),                        //       .clken
		.write2      (onchip_sram_s2_write),                        //       .write
		.readdata2   (onchip_sram_s2_readdata),                     //       .readdata
		.writedata2  (onchip_sram_s2_writedata),                    //       .writedata
		.byteenable2 (onchip_sram_s2_byteenable),                   //       .byteenable
		.clk2        (onchip_sram_clk2_clk),                        //   clk2.clk
		.reset2      (onchip_sram_reset2_reset),                    // reset2.reset
		.reset_req2  (onchip_sram_reset2_reset_req),                //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_dma_1 dma_1 (
		.clk                (system_pll_sys_clk_clk),                                //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                       //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_1_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_1_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_1_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_1_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_1_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (),                                                      //                irq.irq
		.read_address       (dma_1_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_1_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_1_read_master_read),                                //                   .read_n
		.read_readdata      (dma_1_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_1_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_1_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_1_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_1_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_1_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_1_write_master_write),                              //                   .write_n
		.write_writedata    (dma_1_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_1_write_master_byteenable)                          //                   .byteenable
	);

	Computer_System_dma_2 dma_2 (
		.clk                (system_pll_sys_clk_clk),                                //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                       //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_2_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_2_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_2_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_2_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_2_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (),                                                      //                irq.irq
		.read_address       (dma_2_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_2_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_2_read_master_read),                                //                   .read_n
		.read_readdata      (dma_2_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_2_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_2_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_2_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_2_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_2_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_2_write_master_write),                              //                   .write_n
		.write_writedata    (dma_2_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_2_write_master_byteenable)                          //                   .byteenable
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                     //                                       ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                   //                                                                   .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                    //                                                                   .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                   //                                                                   .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                  //                                                                   .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                   //                                                                   .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                  //                                                                   .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                   //                                                                   .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                  //                                                                   .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                  //                                                                   .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                      //                                                                   .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                    //                                                                   .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                    //                                                                   .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                    //                                                                   .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                   //                                                                   .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                   //                                                                   .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                      //                                                                   .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                    //                                                                   .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                   //                                                                   .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                   //                                                                   .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                     //                                                                   .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                   //                                                                   .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                    //                                                                   .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                   //                                                                   .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                  //                                                                   .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                   //                                                                   .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                  //                                                                   .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                   //                                                                   .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                  //                                                                   .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                  //                                                                   .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                      //                                                                   .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                    //                                                                   .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                    //                                                                   .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                    //                                                                   .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                   //                                                                   .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                   //                                                                   .rready
		.System_PLL_sys_clk_clk                                                   (system_pll_sys_clk_clk),                                //                                                 System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // ARM_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.dma_1_reset_reset_bridge_in_reset_reset                                  (rst_controller_reset_out_reset),                        //                                  dma_1_reset_reset_bridge_in_reset.reset
		.dma_1_control_port_slave_address                                         (mm_interconnect_0_dma_1_control_port_slave_address),    //                                           dma_1_control_port_slave.address
		.dma_1_control_port_slave_write                                           (mm_interconnect_0_dma_1_control_port_slave_write),      //                                                                   .write
		.dma_1_control_port_slave_readdata                                        (mm_interconnect_0_dma_1_control_port_slave_readdata),   //                                                                   .readdata
		.dma_1_control_port_slave_writedata                                       (mm_interconnect_0_dma_1_control_port_slave_writedata),  //                                                                   .writedata
		.dma_1_control_port_slave_chipselect                                      (mm_interconnect_0_dma_1_control_port_slave_chipselect), //                                                                   .chipselect
		.dma_2_control_port_slave_address                                         (mm_interconnect_0_dma_2_control_port_slave_address),    //                                           dma_2_control_port_slave.address
		.dma_2_control_port_slave_write                                           (mm_interconnect_0_dma_2_control_port_slave_write),      //                                                                   .write
		.dma_2_control_port_slave_readdata                                        (mm_interconnect_0_dma_2_control_port_slave_readdata),   //                                                                   .readdata
		.dma_2_control_port_slave_writedata                                       (mm_interconnect_0_dma_2_control_port_slave_writedata),  //                                                                   .writedata
		.dma_2_control_port_slave_chipselect                                      (mm_interconnect_0_dma_2_control_port_slave_chipselect)  //                                                                   .chipselect
	);

	Computer_System_mm_interconnect_1 mm_interconnect_1 (
		.ARM_A9_HPS_f2h_axi_slave_awid                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid),    //                                        ARM_A9_HPS_f2h_axi_slave.awid
		.ARM_A9_HPS_f2h_axi_slave_awaddr                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr),  //                                                                .awaddr
		.ARM_A9_HPS_f2h_axi_slave_awlen                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen),   //                                                                .awlen
		.ARM_A9_HPS_f2h_axi_slave_awsize                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize),  //                                                                .awsize
		.ARM_A9_HPS_f2h_axi_slave_awburst                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst), //                                                                .awburst
		.ARM_A9_HPS_f2h_axi_slave_awlock                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock),  //                                                                .awlock
		.ARM_A9_HPS_f2h_axi_slave_awcache                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache), //                                                                .awcache
		.ARM_A9_HPS_f2h_axi_slave_awprot                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot),  //                                                                .awprot
		.ARM_A9_HPS_f2h_axi_slave_awuser                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser),  //                                                                .awuser
		.ARM_A9_HPS_f2h_axi_slave_awvalid                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid), //                                                                .awvalid
		.ARM_A9_HPS_f2h_axi_slave_awready                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready), //                                                                .awready
		.ARM_A9_HPS_f2h_axi_slave_wid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid),     //                                                                .wid
		.ARM_A9_HPS_f2h_axi_slave_wdata                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata),   //                                                                .wdata
		.ARM_A9_HPS_f2h_axi_slave_wstrb                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb),   //                                                                .wstrb
		.ARM_A9_HPS_f2h_axi_slave_wlast                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast),   //                                                                .wlast
		.ARM_A9_HPS_f2h_axi_slave_wvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid),  //                                                                .wvalid
		.ARM_A9_HPS_f2h_axi_slave_wready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready),  //                                                                .wready
		.ARM_A9_HPS_f2h_axi_slave_bid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid),     //                                                                .bid
		.ARM_A9_HPS_f2h_axi_slave_bresp                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp),   //                                                                .bresp
		.ARM_A9_HPS_f2h_axi_slave_bvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid),  //                                                                .bvalid
		.ARM_A9_HPS_f2h_axi_slave_bready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready),  //                                                                .bready
		.ARM_A9_HPS_f2h_axi_slave_arid                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid),    //                                                                .arid
		.ARM_A9_HPS_f2h_axi_slave_araddr                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr),  //                                                                .araddr
		.ARM_A9_HPS_f2h_axi_slave_arlen                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen),   //                                                                .arlen
		.ARM_A9_HPS_f2h_axi_slave_arsize                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize),  //                                                                .arsize
		.ARM_A9_HPS_f2h_axi_slave_arburst                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst), //                                                                .arburst
		.ARM_A9_HPS_f2h_axi_slave_arlock                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock),  //                                                                .arlock
		.ARM_A9_HPS_f2h_axi_slave_arcache                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache), //                                                                .arcache
		.ARM_A9_HPS_f2h_axi_slave_arprot                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot),  //                                                                .arprot
		.ARM_A9_HPS_f2h_axi_slave_aruser                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser),  //                                                                .aruser
		.ARM_A9_HPS_f2h_axi_slave_arvalid                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid), //                                                                .arvalid
		.ARM_A9_HPS_f2h_axi_slave_arready                                      (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready), //                                                                .arready
		.ARM_A9_HPS_f2h_axi_slave_rid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid),     //                                                                .rid
		.ARM_A9_HPS_f2h_axi_slave_rdata                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata),   //                                                                .rdata
		.ARM_A9_HPS_f2h_axi_slave_rresp                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp),   //                                                                .rresp
		.ARM_A9_HPS_f2h_axi_slave_rlast                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast),   //                                                                .rlast
		.ARM_A9_HPS_f2h_axi_slave_rvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid),  //                                                                .rvalid
		.ARM_A9_HPS_f2h_axi_slave_rready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready),  //                                                                .rready
		.System_PLL_sys_clk_clk                                                (system_pll_sys_clk_clk),                             //                                              System_PLL_sys_clk.clk
		.ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                 // ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.dma_1_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),                     //                               dma_1_reset_reset_bridge_in_reset.reset
		.dma_1_read_master_address                                             (dma_1_read_master_address),                          //                                               dma_1_read_master.address
		.dma_1_read_master_waitrequest                                         (dma_1_read_master_waitrequest),                      //                                                                .waitrequest
		.dma_1_read_master_chipselect                                          (dma_1_read_master_chipselect),                       //                                                                .chipselect
		.dma_1_read_master_read                                                (~dma_1_read_master_read),                            //                                                                .read
		.dma_1_read_master_readdata                                            (dma_1_read_master_readdata),                         //                                                                .readdata
		.dma_1_read_master_readdatavalid                                       (dma_1_read_master_readdatavalid),                    //                                                                .readdatavalid
		.dma_2_write_master_address                                            (dma_2_write_master_address),                         //                                              dma_2_write_master.address
		.dma_2_write_master_waitrequest                                        (dma_2_write_master_waitrequest),                     //                                                                .waitrequest
		.dma_2_write_master_byteenable                                         (dma_2_write_master_byteenable),                      //                                                                .byteenable
		.dma_2_write_master_chipselect                                         (dma_2_write_master_chipselect),                      //                                                                .chipselect
		.dma_2_write_master_write                                              (~dma_2_write_master_write),                          //                                                                .write
		.dma_2_write_master_writedata                                          (dma_2_write_master_writedata)                        //                                                                .writedata
	);

	Computer_System_mm_interconnect_2 mm_interconnect_2 (
		.System_PLL_sys_clk_clk                  (system_pll_sys_clk_clk),                      //                System_PLL_sys_clk.clk
		.dma_2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),              // dma_2_reset_reset_bridge_in_reset.reset
		.dma_1_write_master_address              (dma_1_write_master_address),                  //                dma_1_write_master.address
		.dma_1_write_master_waitrequest          (dma_1_write_master_waitrequest),              //                                  .waitrequest
		.dma_1_write_master_byteenable           (dma_1_write_master_byteenable),               //                                  .byteenable
		.dma_1_write_master_chipselect           (dma_1_write_master_chipselect),               //                                  .chipselect
		.dma_1_write_master_write                (~dma_1_write_master_write),                   //                                  .write
		.dma_1_write_master_writedata            (dma_1_write_master_writedata),                //                                  .writedata
		.dma_2_read_master_address               (dma_2_read_master_address),                   //                 dma_2_read_master.address
		.dma_2_read_master_waitrequest           (dma_2_read_master_waitrequest),               //                                  .waitrequest
		.dma_2_read_master_chipselect            (dma_2_read_master_chipselect),                //                                  .chipselect
		.dma_2_read_master_read                  (~dma_2_read_master_read),                     //                                  .read
		.dma_2_read_master_readdata              (dma_2_read_master_readdata),                  //                                  .readdata
		.dma_2_read_master_readdatavalid         (dma_2_read_master_readdatavalid),             //                                  .readdatavalid
		.Onchip_SRAM_s1_address                  (mm_interconnect_2_onchip_sram_s1_address),    //                    Onchip_SRAM_s1.address
		.Onchip_SRAM_s1_write                    (mm_interconnect_2_onchip_sram_s1_write),      //                                  .write
		.Onchip_SRAM_s1_readdata                 (mm_interconnect_2_onchip_sram_s1_readdata),   //                                  .readdata
		.Onchip_SRAM_s1_writedata                (mm_interconnect_2_onchip_sram_s1_writedata),  //                                  .writedata
		.Onchip_SRAM_s1_byteenable               (mm_interconnect_2_onchip_sram_s1_byteenable), //                                  .byteenable
		.Onchip_SRAM_s1_chipselect               (mm_interconnect_2_onchip_sram_s1_chipselect), //                                  .chipselect
		.Onchip_SRAM_s1_clken                    (mm_interconnect_2_onchip_sram_s1_clken)       //                                  .clken
	);

	Computer_System_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
